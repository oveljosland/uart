/* testbench for rx module */