library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.pkg.all;

entity top is
	port ( /* TODO: decide which ports to consider */
		clk: in std_logic; /* SYS_CLK_FRQ defined in pkg */
		rst: in std_logic; /* RST defined in pkg */

		rx: in std_logic; 
		tx: out std_logic;

		seg : out std_logic_vector(6 downto 0)
	);
end entity;

architecture rtl of top is
	signal rx_dv: std_logic;
	signal tx_dv: std_logic;

	signal baud_tick: std_logic;

	/* rx tx io */
	signal rx_dout: std_logic_vector(BITWIDTH - 1 downto 0);
	signal tx_din: std_logic_vector(BITWIDTH - 1 downto 0);
	
	/* rx fifo */
	signal ff_din: std_logic_vector(BITWIDTH - 1 downto 0);
	signal ff_dout: std_logic_vector(BITWIDTH - 1 downto 0);
	signal ff_read, ff_write: std_logic; /* r/w enable */
	signal ff_empty, ff_full: std_logic; /* stauts flags */
begin
	baud_clock: entity work.baud_clock
		port map (
			clk => clk,
			rst => rst,
			baud_tick => baud_tick
		);

	rx_module: entity work.rx
		port map (
			clk => clk,
			rst => rst,
			serial_in => rx,
			baud_tick => baud_tick,
			data_valid => rx_dv,
			byte_out => rx_dout
		);

	rx_fifo: entity work.fifo
		port map (
			clk => clk,
			rst => rst,
			r => ff_read,
			w => rx_dv,
			din => rx_dout,
			dout => ff_dout,
			empty => ff_empty,
			full => ff_full
		);
	display: entity work.display
		port map (
			char => rx_dout,
			seg => seg
		);
end architecture;
