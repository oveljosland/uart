/* testbench for rx module */
/* Denne testbenken skal kunne simulere oppførselen til rx modulen */

