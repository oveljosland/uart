library ieee;
use ieee.std_logic_1164.all;

entity display is
end entity;

architecture rtl of display is
end architecture;